`timescale 1ns / 1ps
module barrelshifter32_tb;
reg [31:0] a;
reg [4:0] b;
reg [1:0] aluc;
wire [31:0] c;
barrelshifter32 uut(
.a(a), 
.b(b), 
.aluc(aluc), 
.c(c));
initial
begin
//������������
a = 32'b00101010010010000010001000010010;
b = 5'b01111;
aluc = 2'b11;
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01010;
aluc = 2'b11;
//�����߼�����
#40
a = 32'b00101010010010000010001000010010;
b = 5'b00100;
aluc = 2'b01;
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01100;
aluc = 2'b01;
//�����߼�����
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01010;
aluc = 2'b10;
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01010;
aluc = 2'b10;
//������������
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01010;
aluc = 2'b00;
#40
a = 32'b00101010010010000010001000010010;
b = 5'b01010;
aluc = 2'b00;
end
endmodule